`timescale 1 ns / 100 ps
package STATES;
    typedef enum reg [1:0] {FETCH, DECODE, EXECUTE, UPDATE} PHASES;
endpackage
